* MOSFET amplifier
.subckt mosfet g s d
Cgs g s cgs
Gm s d g s gm
Ro d s ro
.end

R0 vin vinx Rs
X0 mosfet vinx 0 vout

P1 vin 0
P2 vout 0

.print Z(1, 1)
.print Y(1, 1)
.print Z(2, 2)
.print Y(2, 2)
