V0 vin 0 1
R1 vin vout 1000
R2 vout 0 1000

.print V(vout)
