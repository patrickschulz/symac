RR1 vin vout R1
RR2 vout 0 R2
VV0 vin 0 V0

*.print V(vout)
*.print I(R1)

.print all
