R0 vx 0 R0
C0 vx 0 C0
