R1 in out foo

.subckt mosfet g d s
R0 p n R0
.end

O2 1 2 3
