.subckt mosfet g s d
C g s cgs
G s d g s gm
R d s ro
.end

.subckt sub p n
R p n R0
.end

V vin 0 vin
Xsub vin 0
