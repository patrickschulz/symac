*Test for subckts
