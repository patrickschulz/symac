Title
R 1 0 R1
* empty line

* second title
Second Title
* wrong component
R 1 2 3 R0
