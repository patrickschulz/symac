* comment
R 1 2 foo
O 1 2 3 bar
.print V(out)
