* Mapping Test
V A 0 V0
R A 0 R0
