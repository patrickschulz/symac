.print 2.5
