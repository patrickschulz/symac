V A 0 Vin
R A B R1
C B 0 C1
