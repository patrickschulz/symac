Vin 1 0 V1
C1 1 2 C1
R1 2 3 R1
C2 3 0 C2    
