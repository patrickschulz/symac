V0 in 0 Vin
V0 in 0 Vin

R1 in out R1

.print V(vout)
