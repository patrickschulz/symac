R1 v1 v1cp z11
F1 v1cn 0 v2cp v2cn z12
R2 v2 v2cp z22
F2 v2cn 0 v1cp v1cn z21

P1 v1 0
P2 v2 0
