* Mapping Test
V A 0 V0
C A 0 R0
