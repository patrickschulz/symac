* MOSFET amplifier
.subckt mosfet g s d
Ggm s d g s gm
Rro d s ro
.end

V0 vin 0 vin
*X1 mosfet vin 0 vout
X mosfet vout 0 vout

*.print all
*.print V(vout)
