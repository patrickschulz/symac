Title
R0 1 0 R1
* empty line

* second title
Second Title
* wrong component
R0 1 2 3 R0
