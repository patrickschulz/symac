* CCVS test
V0 vin 0 Vin
Rin vin vx Rin
Rout vout 0 Rout
F0 vout 0 vx 0 Rtrans

.print I(V0.n)
.print I(F0.cp)
.print I(Rout.p)
.print I(F0.p)
