.subckt mosfet g d s
G s d g s gm
R d s ro
.end

V vin 0 vin
Xmosfet vin vout 0

result print v(vout)
