* MOSFET amplifier
.subckt mosfet g s d
Cgs g s cgs
Gm s d g s gm
Ro d s ro
.end

X0 mosfet vin 0 vout

P1 vin 0
P2 vout 0

.print H(1, 1)
.print H(1, 2)
.print H(2, 1)
.print H(2, 2)
*.print G(1, 1)
*.print G(1, 2)
*.print G(2, 1)
*.print G(2, 2)
