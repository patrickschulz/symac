* MOSFET amplifier
.subckt mosfet g s d
Ccgs g s cgs
Ggm s d g s gm
Rro d s ro
.end

VV0 vinx 0 vin
RV0 vinx vin Rs
X0 mosfet vin 0 vout

.print V(vout)
