Transfer function
V vin 0 Vin
R vin vout R0
R vout 0 R1
