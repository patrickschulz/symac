R1 v1 0 R1
R2 v1 v2 R2

P1 v1 0
P2 v2 0
