* MOSFET amplifier
.subckt mosfet g s d
Cgs g s cgs
Gm s d g s gm
Ro d s ro
.end

V0 vin 0 vin
R0 vin vinx Rs
X0 mosfet vinx 0 vout

.print V(vout) / V(vin)
