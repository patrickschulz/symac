- Voltage sources test
V 1 0 V1
R 1 0 R1
V 2 0 V2
R 2 0 R2
