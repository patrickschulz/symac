Transfer function
V vin 0 Vin
C vout 0 C1
R vin vout R1
