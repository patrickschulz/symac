.command simplify
level english
R1 >> R2 
C1 >> C2
.end

V in 0 Vin
R in 1 R1
C 1 0  C1
R 1 out R2
C out 0 C2
