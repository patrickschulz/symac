* Transistors terminals in the following order: gate drain source
*MP1 vbias vout vdd
*MN1 vin vout vss
*
*Vdd vdd 0 vdd
*Vss vss 0 0
*Vin vin 0 vin

* simpler example: resistance with voltage source
R0 vdd vout RL
M0 vin vout 0
V0 vdd 0 vdd 

.print I(R0.p)
