* Voltage controlled voltage source
VV0 vin 0 vin
RR0 vout 0 Ro
GG0 0 vout vin 0 gm

.print V(vout)
.print I(R0.p)
