I0 vin 0 iin

R0 vin 0 { R0 * A0 }

.print V(vin)
