- CCVS test
R 1 2 Rin
R 3 0 Rout
V 1 0 Vin
H 0 3 2 0 gain
