V 1 0 V0
R 1 2 R1
R 2 0 R2
