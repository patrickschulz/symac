R0 vin vout
