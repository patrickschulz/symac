* MOSFET amplifier
.subckt mosfet g s d
Cgs g s cgs
Gm s d g s gm
Ro d s ro
.end

V0 vinx 0 vin
R0 vinx vin Rs
X0 mosfet vin 0 vout

.print V(vout)
