simulator lang=spectre

R0 in out R0
G0 1 2 3 4 gm
O0 1 2 3

* comment with several words
// spectre-type comment
