- Lowpass
V0 vin 0 vin
R0 vin vout R
C0 vout 0 C

.print V(vout)
