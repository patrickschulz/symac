*Einfacher Mosfet ( ohne Kapazitäten)
.subckt mosfet g s d
.