- MOSFET amplifier
V 1 0 Vin
G 0 2 1 0 gm
R 2 0 Rout
C 2 0 Cout
C 1 3 Cff
R 3 2 Rff
