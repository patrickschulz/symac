R0 vx 0 R0
R1 vx 0 R1
C0 vx 0 C0

.print VN(vx)
