.subckt sub p n
R1 p !out R1
R2 !out n R2
R3 p !0 R3
.end

V0 vin 0 vin
Xsub sub vin 0

*.print all
.print V(!out)
