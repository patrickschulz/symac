R1 v1x v1c h11
E1 v1c 0 v2 0 h12
R2 v2 0 {1/h22}
H2 0 v2 v1 v1x h21

P1 v1 0
P2 v2 0

.print H(1, 1)
.print H(1, 2)
.print H(2, 1)
.print H(2, 2)
