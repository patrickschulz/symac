V0 vout 0 vout
R0 vout 0 Rout

.print I(R0.p)
.print I(R0.n)
