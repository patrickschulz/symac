Transfer function
V vin 0 Vin
R vin 0 R0
