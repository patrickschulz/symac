Transfer function
V vin 0 Vin
R vin vout R1
R vout 0 R2
