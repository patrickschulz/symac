.subckt sub p n
* comment
R2 p n R2
.end

V0 vin 0 vin
X sub vin 0

.print all
