- Subcircuits
.subckt amplifier 
