I 1 0 I0
R 1 0 R0
