R in out R0
G 1 2 3 4 gm
O 1 2 3

* comment with several words
