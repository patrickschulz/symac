* CCVS test
V vin 0 Vin
R vin vx Rin
R vout 0 Rout
F vout 0 vx 0 Rtrans

.print V(vx)
.print V(vout)
