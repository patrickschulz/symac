* Numeric Test
VV0 vin 0 1
RR1 vin vout 1000
RR2 vout 0 1000

.print V(vout)
