R1 v1 v2 Z

P1 v1 0
P2 v2 0

.print ABCD(1, 1)
.print ABCD(1, 2)
.print ABCD(2, 1)
.print ABCD(2, 2)
