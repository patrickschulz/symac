* Voltage controlled current source
V0 vin 0 vin
R0 vout 0 Ro
G0 0 vout vin 0 gm

.print V(vout)
.print I(R0.p)
