Gm1 0 vs vin 0 gm
Rout1 vs 0 rout
Gm2 vs vout vbias vs gm
Rout2 vout vs rout

* capacitances
Cl vout 0 Cl
Cs vs 0 Cs

Vbias vbias 0 0
Vin vin 0 vin

.print V(vout) / V(vin)
