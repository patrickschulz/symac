* Opamp inverter
V0 vin 0 Vin
Rf vin vx Rf
Rfb vx vout Rfb
Op 0 vx vout

.print V(vout) / V(vin)
