- MOSFET amplifier
.subckt mosfet g s d
Cgs g s cgs
G s d g s gm
Ro d s ro
.end

V0 vin 0 vin
X1 mosfet vin 0 vout
Rl vout 0 ro

.print V(vout)
.print all
