.subckt sub p n out
R1 p out R1
R2 out n R2
.end

V0 vin 0 vin
Xsub sub vin 0 vout

*.print all
.print V(vin) / V(vout)
.print V(vin)
