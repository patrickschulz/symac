- Numeric Test
I 1 0 1
R 1 0 50
