* Numeric Test
I0 vout 0 1
R0 vout 0 50

.print V(vout)
