R 1 2 foo
