R0 v1 0 R0

P0 v1 0
