* CCVS test
V0 vin 0 Vin
R1 vin vx Rin
R2 vout 0 Rout
H0 0 vout vx 0 gain

.print V(vx)
.print V(vout)
