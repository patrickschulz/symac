V 1 0 Vin
O 1 2 3
R 3 2 R1
R 2 0 R2
