Mp vbias vout vdd
Mn vin vout 0
Vdd vdd 0 vdd 
Vbias vbias 0 vbias
Vin vin 0 vin ac=1

.print V(vout) / V(vin)
