- Naming Nodes
V vin 0 V1
R vin 0 R1
