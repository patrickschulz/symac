R1 v1 0 R1
R2 v1 v2 R2

P1 v1 0
P2 v2 0

*V1 v1 0 v1
*V2 v2 0 0
*.print -I(V1.p) / V(v1)
*.print -I(V2.p) / V(v1)
