R1 v1 0 1/y11
G1 0 v1 v2 0 y12
R2 v2 0 1/y22
G2 0 v2 v1 0 y21

P1 v1 0
P2 v2 0
