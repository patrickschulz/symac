- MOSFET amplifier
V 1 0 Vin
R 1 2 Rs
C 2 0 Cgs
G 0 3 2 0 gm
R 3 0 Rout
C 3 0 Cout
C 2 4 Cff
R 4 3 Rff
