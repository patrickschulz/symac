- CCVS test
R 1 2 Rin
R 3 0 Rout
V 1 0 Vin
F 3 0 2 0 Rtrans
