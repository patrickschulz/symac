R vin vout R1
R vout 0 R2
V vin 0 V0

*.print V(vout)
*.print I(R1)

.print all
