Gm 0 vout vin 0 gm
Rout vout 0 rout
Cout vout 0 cout

V0 vin 0 vin

In vout 0 0 noise=In

.print VN(vout)
.print VNI(vout)
