*R0 v1 0 R0
R1 v1 vx R1
R2 vx 0 R2

P0 v1 0
*V0 v1 0 v0
