simulator lang=spectre
R0 (in out) resistor R0

simulator lang=spice
V0 in 0 Vin
C0 out 0 Cl

* comment with several words
// spectre-type comment

.print V(out)
